`ifndef CYCLE
    `define CYCLE 10 
`endif //__CYCLE_H___
`timescale 1ns/1ns
