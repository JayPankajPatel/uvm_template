`ifndef __TB_VEND___ // make sure the files are included only once
`define __TB_VEND___ 
    `include "uvm_macros.svh"
    package tb_pkg;
        import uvm_pkg::*; 
    endpackage : tb_pkg

`endif // __TB_VEND___
