module tb_top(); 
    import uvm_pkg::*; 
    import tb_pkg::*; 
    initial begin 
        run_test("test"); 
    end
endmodule : tb_top
